*--------------------------------------
* BAND-PASS ACTIVE FILTER 			  -
*                                     -
* Author: Van Dessel Stijn            -
* Date: 9 may 2018                    -
* Filename: AFtrap_21_mcr5_tl084.cir -
*--------------------------------------
.inc TL084.cir

.model rmod  res(r = 1k  DEV  5%)
.model cmod  cap(c = 1n  DEV 20%)

Vin 7 0 AC 1V
Vcc 10 0  DC  15V
Vee 20 0  DC -15V

R1 5 7 rmod 7.9577
R2 2 3 rmod 7.9577
R3 3 4 rmod 7.9577
R4 4 5 rmod 7.9577
R5 5 6 rmod 15.915
R6 1 6 rmod 7.9577
C1 1 2 cmod 10
C2 5 6 cmod 40

*       i+ i- V+ V-  O
XTL084_1   0  3 10 20  2 TL084
XTL084_2   0  5 10 20  6 TL084
XTL084_3   1  0 10 20  4 TL084

.AC DEC 100 100HZ 10KHZ
.MC 10 AC V(6) YMAX LIST OUTPUT ALL

.PROBE
.END
